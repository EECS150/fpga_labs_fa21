module nco(
    input clk,
    input rst,
    input [23:0] fcw,
    output [9:0] out
);
    assign out = 0;
endmodule
